
/**
 * A mapping from instruction opcodes to mnemonics for instruction tracing during simulation.
 * This module is not used during synthesis.
 */
module Instructions();
    reg [32:0] instruction_map[0:255];
    initial begin
        instruction_map[0] = "HLT ";
        instruction_map[1] = "NOP ";
        instruction_map[2] = "SF  ";
        instruction_map[3] = "RF  ";
        instruction_map[4] = "EI  ";
        instruction_map[5] = "DI  ";
        instruction_map[6] = "SL  ";
        instruction_map[7] = "RL  ";
        instruction_map[8] = "CL  ";
        instruction_map[9] = "RSR ";
        instruction_map[10] = "RI  ";
        instruction_map[11] = "RIM ";
        instruction_map[12] = "ELO ";
        instruction_map[13] = "PCX ";
        instruction_map[14] = "DLY ";
        instruction_map[15] = "RSYS";
        instruction_map[16] = "BL  ";
        instruction_map[17] = "BNL ";
        instruction_map[18] = "BF  ";
        instruction_map[19] = "BNF ";
        instruction_map[20] = "BZ  ";
        instruction_map[21] = "BNZ ";
        instruction_map[22] = "BM  ";
        instruction_map[23] = "BP  ";
        instruction_map[24] = "BGZ ";
        instruction_map[25] = "BLE ";
        instruction_map[26] = "BS1 ";
        instruction_map[27] = "BS2 ";
        instruction_map[28] = "BS3 ";
        instruction_map[29] = "BS4 ";
        instruction_map[30] = "BTM?";
        instruction_map[31] = "BEP?";
        instruction_map[32] = "INR ";
        instruction_map[33] = "DCR ";
        instruction_map[34] = "CLR ";
        instruction_map[35] = "IVR ";
        instruction_map[36] = "SRR ";
        instruction_map[37] = "SLR ";
        instruction_map[38] = "RRR ";
        instruction_map[39] = "RLR ";
        instruction_map[40] = "INAL";
        instruction_map[41] = "DCAL";
        instruction_map[42] = "CLAL";
        instruction_map[43] = "IVAL";
        instruction_map[44] = "SRAL";
        instruction_map[45] = "SLAL";
        instruction_map[46] = "?2e ";
        instruction_map[47] = "?2f ";
        instruction_map[48] = "INRW";
        instruction_map[49] = "DCR ";
        instruction_map[50] = "CLR ";
        instruction_map[51] = "IVR ";
        instruction_map[52] = "SRR ";
        instruction_map[53] = "SLR ";
        instruction_map[54] = "RRR ";
        instruction_map[55] = "RLR ";
        instruction_map[56] = "INAW";
        instruction_map[57] = "DCAW";
        instruction_map[58] = "CLAW";
        instruction_map[59] = "IVAW";
        instruction_map[60] = "SRAW";
        instruction_map[61] = "SLAW";
        instruction_map[62] = "INX ";
        instruction_map[63] = "DCX ";
        instruction_map[64] = "ADD ";
        instruction_map[65] = "SUB ";
        instruction_map[66] = "AND ";
        instruction_map[67] = "ORI ";
        instruction_map[68] = "ORE ";
        instruction_map[69] = "XFR ";
        instruction_map[70] = "?46 ";
        instruction_map[71] = "?47 ";
        instruction_map[72] = "AABL";
        instruction_map[73] = "SABL";
        instruction_map[74] = "NABL";
        instruction_map[75] = "XAXL";
        instruction_map[76] = "XAYL";
        instruction_map[77] = "XABL";
        instruction_map[78] = "XAZL";
        instruction_map[79] = "XASL";
        instruction_map[80] = "ADD ";
        instruction_map[81] = "SUB ";
        instruction_map[82] = "AND ";
        instruction_map[83] = "ORI ";
        instruction_map[84] = "ORE ";
        instruction_map[85] = "XFR ";
        instruction_map[86] = "?56 ";
        instruction_map[87] = "?57 ";
        instruction_map[88] = "AABW";
        instruction_map[89] = "SABW";
        instruction_map[90] = "NABW";
        instruction_map[91] = "XAXW";
        instruction_map[92] = "XAYW";
        instruction_map[93] = "XABW";
        instruction_map[94] = "XAZW";
        instruction_map[95] = "XASW";
        instruction_map[96] = "LDXW";
        instruction_map[97] = "LDXW";
        instruction_map[98] = "LDXW";
        instruction_map[99] = "LDXW";
        instruction_map[100] = "LDXW";
        instruction_map[101] = "LDXW";
        instruction_map[102] = "JSYS";
        instruction_map[103] = "?67 ";
        instruction_map[104] = "STXW";
        instruction_map[105] = "STXW";
        instruction_map[106] = "STXW";
        instruction_map[107] = "STXW";
        instruction_map[108] = "STXW";
        instruction_map[109] = "STXW";
        instruction_map[110] = "LDCC";
        instruction_map[111] = "STCC";
        instruction_map[112] = "JMP ";
        instruction_map[113] = "JMP ";
        instruction_map[114] = "JMP ";
        instruction_map[115] = "JMP ";
        instruction_map[116] = "JMP ";
        instruction_map[117] = "JMP ";
        instruction_map[118] = "?76 ";
        instruction_map[119] = "?77 ";
        instruction_map[120] = "?78 ";
        instruction_map[121] = "JSR ";
        instruction_map[122] = "JSR ";
        instruction_map[123] = "JSR ";
        instruction_map[124] = "JSR ";
        instruction_map[125] = "JSR ";
        instruction_map[126] = "PUSH";
        instruction_map[127] = "POP ";
        instruction_map[128] = "LDAL";
        instruction_map[129] = "LDAL";
        instruction_map[130] = "LDAL";
        instruction_map[131] = "LDAL";
        instruction_map[132] = "LDAL";
        instruction_map[133] = "LDAL";
        instruction_map[134] = "?86 ";
        instruction_map[135] = "?87 ";
        instruction_map[136] = "LALA";
        instruction_map[137] = "LALB";
        instruction_map[138] = "LALX";
        instruction_map[139] = "LALY";
        instruction_map[140] = "LALZ";
        instruction_map[141] = "LALS";
        instruction_map[142] = "LALC";
        instruction_map[143] = "LALP";
        instruction_map[144] = "LDAW";
        instruction_map[145] = "LDAW";
        instruction_map[146] = "LDAW";
        instruction_map[147] = "LDAW";
        instruction_map[148] = "LDAW";
        instruction_map[149] = "LDAW";
        instruction_map[150] = "?96 ";
        instruction_map[151] = "?97 ";
        instruction_map[152] = "LAWA";
        instruction_map[153] = "LAWB";
        instruction_map[154] = "LAWX";
        instruction_map[155] = "LAWY";
        instruction_map[156] = "LAWZ";
        instruction_map[157] = "LAWS";
        instruction_map[158] = "LAWC";
        instruction_map[159] = "LAWP";
        instruction_map[160] = "STAL";
        instruction_map[161] = "STAL";
        instruction_map[162] = "STAL";
        instruction_map[163] = "STAL";
        instruction_map[164] = "STAL";
        instruction_map[165] = "STAL";
        instruction_map[166] = "?a6 ";
        instruction_map[167] = "?a7 ";
        instruction_map[168] = "SALA";
        instruction_map[169] = "SALB";
        instruction_map[170] = "SALX";
        instruction_map[171] = "SALY";
        instruction_map[172] = "SALZ";
        instruction_map[173] = "SALS";
        instruction_map[174] = "SALC";
        instruction_map[175] = "SALP";
        instruction_map[176] = "STAW";
        instruction_map[177] = "STAW";
        instruction_map[178] = "STAW";
        instruction_map[179] = "STAW";
        instruction_map[180] = "STAW";
        instruction_map[181] = "STAW";
        instruction_map[182] = "?b6 ";
        instruction_map[183] = "?b7 ";
        instruction_map[184] = "SAWA";
        instruction_map[185] = "SAWB";
        instruction_map[186] = "SAWX";
        instruction_map[187] = "SAWY";
        instruction_map[188] = "SAWZ";
        instruction_map[189] = "SAWS";
        instruction_map[190] = "SAWC";
        instruction_map[191] = "SAWP";
        instruction_map[192] = "LDBL";
        instruction_map[193] = "LDBL";
        instruction_map[194] = "LDBL";
        instruction_map[195] = "LDBL";
        instruction_map[196] = "LDBL";
        instruction_map[197] = "LDBL";
        instruction_map[198] = "?c6 ";
        instruction_map[199] = "?c7 ";
        instruction_map[200] = "LBLA";
        instruction_map[201] = "LBLB";
        instruction_map[202] = "LBLX";
        instruction_map[203] = "LBLY";
        instruction_map[204] = "LBLZ";
        instruction_map[205] = "LBLS";
        instruction_map[206] = "LBLC";
        instruction_map[207] = "LBLP";
        instruction_map[208] = "LDBW";
        instruction_map[209] = "LDBW";
        instruction_map[210] = "LDBW";
        instruction_map[211] = "LDBW";
        instruction_map[212] = "LDBW";
        instruction_map[213] = "LDBW";
        instruction_map[214] = "?d6 ";
        instruction_map[215] = "?d7 ";
        instruction_map[216] = "LBWA";
        instruction_map[217] = "LBWB";
        instruction_map[218] = "LBWX";
        instruction_map[219] = "LDBW";
        instruction_map[220] = "LBWZ";
        instruction_map[221] = "LBWS";
        instruction_map[222] = "LBWC";
        instruction_map[223] = "LBWP";
        instruction_map[224] = "STBL";
        instruction_map[225] = "STBL";
        instruction_map[226] = "STBL";
        instruction_map[227] = "STBL";
        instruction_map[228] = "STBL";
        instruction_map[229] = "STBL";
        instruction_map[230] = "?e6 ";
        instruction_map[231] = "?e7 ";
        instruction_map[232] = "SBLA";
        instruction_map[233] = "SBLB";
        instruction_map[234] = "SBLX";
        instruction_map[235] = "SBLY";
        instruction_map[236] = "SBLZ";
        instruction_map[237] = "SBLS";
        instruction_map[238] = "SBLC";
        instruction_map[239] = "SBLP";
        instruction_map[240] = "STBW";
        instruction_map[241] = "STBW";
        instruction_map[242] = "STBW";
        instruction_map[243] = "STBW";
        instruction_map[244] = "STBW";
        instruction_map[245] = "STBW";
        instruction_map[246] = "?f6 ";
        instruction_map[247] = "?f7 ";
        instruction_map[248] = "SBWA";
        instruction_map[249] = "SBWB";
        instruction_map[250] = "SBWX";
        instruction_map[251] = "SBWY";
        instruction_map[252] = "SBWZ";
        instruction_map[253] = "SBWS";
        instruction_map[254] = "SBWC";
        instruction_map[255] = "SBWP";
    end
endmodule
